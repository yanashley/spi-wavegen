module top(
    input logic     clk,
    input logic     rst,

    // output logics will be same as MP3 prob
);
endmodule
